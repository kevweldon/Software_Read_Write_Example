module sys (
		input  wire       clk_clk,         //      clk.clk
		output wire [7:0] pio_8bit_export, // pio_8bit.export
		input  wire       reset_reset      //    reset.reset
	);
endmodule

