// sys.v

// Generated using ACDS version 21.4 67

`timescale 1 ps / 1 ps
module sys (
		input  wire       clk_clk,         //      clk.clk
		output wire [7:0] pio_8bit_export, // pio_8bit.export
		input  wire       reset_reset      //    reset.reset
	);

	wire         clock_in_out_clk_clk;                                      // clock_in:out_clk -> [cpu:clk, data_instruction_ram:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:clock_in_out_clk_clk, pio_8bit:clk, ram_32bit:clk, reset_in:clk, rst_controller:clk]
	wire  [31:0] cpu_data_manager_awaddr;                                   // cpu:data_manager_awaddr -> mm_interconnect_0:cpu_data_manager_awaddr
	wire   [1:0] cpu_data_manager_bresp;                                    // mm_interconnect_0:cpu_data_manager_bresp -> cpu:data_manager_bresp
	wire         cpu_data_manager_arready;                                  // mm_interconnect_0:cpu_data_manager_arready -> cpu:data_manager_arready
	wire  [31:0] cpu_data_manager_rdata;                                    // mm_interconnect_0:cpu_data_manager_rdata -> cpu:data_manager_rdata
	wire   [3:0] cpu_data_manager_wstrb;                                    // cpu:data_manager_wstrb -> mm_interconnect_0:cpu_data_manager_wstrb
	wire         cpu_data_manager_wready;                                   // mm_interconnect_0:cpu_data_manager_wready -> cpu:data_manager_wready
	wire         cpu_data_manager_awready;                                  // mm_interconnect_0:cpu_data_manager_awready -> cpu:data_manager_awready
	wire         cpu_data_manager_rready;                                   // cpu:data_manager_rready -> mm_interconnect_0:cpu_data_manager_rready
	wire   [2:0] cpu_data_manager_arsize;                                   // cpu:data_manager_arsize -> mm_interconnect_0:cpu_data_manager_arsize
	wire         cpu_data_manager_bready;                                   // cpu:data_manager_bready -> mm_interconnect_0:cpu_data_manager_bready
	wire         cpu_data_manager_wlast;                                    // cpu:data_manager_wlast -> mm_interconnect_0:cpu_data_manager_wlast
	wire         cpu_data_manager_wvalid;                                   // cpu:data_manager_wvalid -> mm_interconnect_0:cpu_data_manager_wvalid
	wire  [31:0] cpu_data_manager_araddr;                                   // cpu:data_manager_araddr -> mm_interconnect_0:cpu_data_manager_araddr
	wire   [2:0] cpu_data_manager_arprot;                                   // cpu:data_manager_arprot -> mm_interconnect_0:cpu_data_manager_arprot
	wire   [1:0] cpu_data_manager_rresp;                                    // mm_interconnect_0:cpu_data_manager_rresp -> cpu:data_manager_rresp
	wire   [2:0] cpu_data_manager_awprot;                                   // cpu:data_manager_awprot -> mm_interconnect_0:cpu_data_manager_awprot
	wire  [31:0] cpu_data_manager_wdata;                                    // cpu:data_manager_wdata -> mm_interconnect_0:cpu_data_manager_wdata
	wire         cpu_data_manager_arvalid;                                  // cpu:data_manager_arvalid -> mm_interconnect_0:cpu_data_manager_arvalid
	wire         cpu_data_manager_bvalid;                                   // mm_interconnect_0:cpu_data_manager_bvalid -> cpu:data_manager_bvalid
	wire   [2:0] cpu_data_manager_awsize;                                   // cpu:data_manager_awsize -> mm_interconnect_0:cpu_data_manager_awsize
	wire         cpu_data_manager_awvalid;                                  // cpu:data_manager_awvalid -> mm_interconnect_0:cpu_data_manager_awvalid
	wire         cpu_data_manager_rvalid;                                   // mm_interconnect_0:cpu_data_manager_rvalid -> cpu:data_manager_rvalid
	wire  [31:0] cpu_instruction_manager_awaddr;                            // cpu:instruction_manager_awaddr -> mm_interconnect_0:cpu_instruction_manager_awaddr
	wire   [1:0] cpu_instruction_manager_bresp;                             // mm_interconnect_0:cpu_instruction_manager_bresp -> cpu:instruction_manager_bresp
	wire         cpu_instruction_manager_arready;                           // mm_interconnect_0:cpu_instruction_manager_arready -> cpu:instruction_manager_arready
	wire  [31:0] cpu_instruction_manager_rdata;                             // mm_interconnect_0:cpu_instruction_manager_rdata -> cpu:instruction_manager_rdata
	wire   [3:0] cpu_instruction_manager_wstrb;                             // cpu:instruction_manager_wstrb -> mm_interconnect_0:cpu_instruction_manager_wstrb
	wire         cpu_instruction_manager_wready;                            // mm_interconnect_0:cpu_instruction_manager_wready -> cpu:instruction_manager_wready
	wire         cpu_instruction_manager_awready;                           // mm_interconnect_0:cpu_instruction_manager_awready -> cpu:instruction_manager_awready
	wire         cpu_instruction_manager_rready;                            // cpu:instruction_manager_rready -> mm_interconnect_0:cpu_instruction_manager_rready
	wire   [2:0] cpu_instruction_manager_arsize;                            // cpu:instruction_manager_arsize -> mm_interconnect_0:cpu_instruction_manager_arsize
	wire         cpu_instruction_manager_bready;                            // cpu:instruction_manager_bready -> mm_interconnect_0:cpu_instruction_manager_bready
	wire         cpu_instruction_manager_wlast;                             // cpu:instruction_manager_wlast -> mm_interconnect_0:cpu_instruction_manager_wlast
	wire         cpu_instruction_manager_wvalid;                            // cpu:instruction_manager_wvalid -> mm_interconnect_0:cpu_instruction_manager_wvalid
	wire  [31:0] cpu_instruction_manager_araddr;                            // cpu:instruction_manager_araddr -> mm_interconnect_0:cpu_instruction_manager_araddr
	wire   [2:0] cpu_instruction_manager_arprot;                            // cpu:instruction_manager_arprot -> mm_interconnect_0:cpu_instruction_manager_arprot
	wire   [1:0] cpu_instruction_manager_rresp;                             // mm_interconnect_0:cpu_instruction_manager_rresp -> cpu:instruction_manager_rresp
	wire   [2:0] cpu_instruction_manager_awprot;                            // cpu:instruction_manager_awprot -> mm_interconnect_0:cpu_instruction_manager_awprot
	wire  [31:0] cpu_instruction_manager_wdata;                             // cpu:instruction_manager_wdata -> mm_interconnect_0:cpu_instruction_manager_wdata
	wire         cpu_instruction_manager_arvalid;                           // cpu:instruction_manager_arvalid -> mm_interconnect_0:cpu_instruction_manager_arvalid
	wire         cpu_instruction_manager_bvalid;                            // mm_interconnect_0:cpu_instruction_manager_bvalid -> cpu:instruction_manager_bvalid
	wire   [2:0] cpu_instruction_manager_awsize;                            // cpu:instruction_manager_awsize -> mm_interconnect_0:cpu_instruction_manager_awsize
	wire         cpu_instruction_manager_awvalid;                           // cpu:instruction_manager_awvalid -> mm_interconnect_0:cpu_instruction_manager_awvalid
	wire         cpu_instruction_manager_rvalid;                            // mm_interconnect_0:cpu_instruction_manager_rvalid -> cpu:instruction_manager_rvalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_dm_agent_readdata;                   // cpu:dm_agent_readdata -> mm_interconnect_0:cpu_dm_agent_readdata
	wire         mm_interconnect_0_cpu_dm_agent_waitrequest;                // cpu:dm_agent_waitrequest -> mm_interconnect_0:cpu_dm_agent_waitrequest
	wire  [15:0] mm_interconnect_0_cpu_dm_agent_address;                    // mm_interconnect_0:cpu_dm_agent_address -> cpu:dm_agent_address
	wire         mm_interconnect_0_cpu_dm_agent_read;                       // mm_interconnect_0:cpu_dm_agent_read -> cpu:dm_agent_read
	wire         mm_interconnect_0_cpu_dm_agent_readdatavalid;              // cpu:dm_agent_readdatavalid -> mm_interconnect_0:cpu_dm_agent_readdatavalid
	wire         mm_interconnect_0_cpu_dm_agent_write;                      // mm_interconnect_0:cpu_dm_agent_write -> cpu:dm_agent_write
	wire  [31:0] mm_interconnect_0_cpu_dm_agent_writedata;                  // mm_interconnect_0:cpu_dm_agent_writedata -> cpu:dm_agent_writedata
	wire         mm_interconnect_0_data_instruction_ram_s1_chipselect;      // mm_interconnect_0:data_instruction_ram_s1_chipselect -> data_instruction_ram:chipselect
	wire  [31:0] mm_interconnect_0_data_instruction_ram_s1_readdata;        // data_instruction_ram:readdata -> mm_interconnect_0:data_instruction_ram_s1_readdata
	wire  [16:0] mm_interconnect_0_data_instruction_ram_s1_address;         // mm_interconnect_0:data_instruction_ram_s1_address -> data_instruction_ram:address
	wire   [3:0] mm_interconnect_0_data_instruction_ram_s1_byteenable;      // mm_interconnect_0:data_instruction_ram_s1_byteenable -> data_instruction_ram:byteenable
	wire         mm_interconnect_0_data_instruction_ram_s1_write;           // mm_interconnect_0:data_instruction_ram_s1_write -> data_instruction_ram:write
	wire  [31:0] mm_interconnect_0_data_instruction_ram_s1_writedata;       // mm_interconnect_0:data_instruction_ram_s1_writedata -> data_instruction_ram:writedata
	wire         mm_interconnect_0_data_instruction_ram_s1_clken;           // mm_interconnect_0:data_instruction_ram_s1_clken -> data_instruction_ram:clken
	wire         mm_interconnect_0_ram_32bit_s1_chipselect;                 // mm_interconnect_0:ram_32bit_s1_chipselect -> ram_32bit:chipselect
	wire  [31:0] mm_interconnect_0_ram_32bit_s1_readdata;                   // ram_32bit:readdata -> mm_interconnect_0:ram_32bit_s1_readdata
	wire   [5:0] mm_interconnect_0_ram_32bit_s1_address;                    // mm_interconnect_0:ram_32bit_s1_address -> ram_32bit:address
	wire   [3:0] mm_interconnect_0_ram_32bit_s1_byteenable;                 // mm_interconnect_0:ram_32bit_s1_byteenable -> ram_32bit:byteenable
	wire         mm_interconnect_0_ram_32bit_s1_write;                      // mm_interconnect_0:ram_32bit_s1_write -> ram_32bit:write
	wire  [31:0] mm_interconnect_0_ram_32bit_s1_writedata;                  // mm_interconnect_0:ram_32bit_s1_writedata -> ram_32bit:writedata
	wire         mm_interconnect_0_ram_32bit_s1_clken;                      // mm_interconnect_0:ram_32bit_s1_clken -> ram_32bit:clken
	wire         mm_interconnect_0_pio_8bit_s1_chipselect;                  // mm_interconnect_0:pio_8bit_s1_chipselect -> pio_8bit:chipselect
	wire  [31:0] mm_interconnect_0_pio_8bit_s1_readdata;                    // pio_8bit:readdata -> mm_interconnect_0:pio_8bit_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_8bit_s1_address;                     // mm_interconnect_0:pio_8bit_s1_address -> pio_8bit:address
	wire         mm_interconnect_0_pio_8bit_s1_write;                       // mm_interconnect_0:pio_8bit_s1_write -> pio_8bit:write_n
	wire  [31:0] mm_interconnect_0_pio_8bit_s1_writedata;                   // mm_interconnect_0:pio_8bit_s1_writedata -> pio_8bit:writedata
	wire  [31:0] mm_interconnect_0_cpu_timer_sw_agent_readdata;             // cpu:timer_sw_agent_readdata -> mm_interconnect_0:cpu_timer_sw_agent_readdata
	wire   [5:0] mm_interconnect_0_cpu_timer_sw_agent_address;              // mm_interconnect_0:cpu_timer_sw_agent_address -> cpu:timer_sw_agent_address
	wire         mm_interconnect_0_cpu_timer_sw_agent_read;                 // mm_interconnect_0:cpu_timer_sw_agent_read -> cpu:timer_sw_agent_read
	wire   [3:0] mm_interconnect_0_cpu_timer_sw_agent_byteenable;           // mm_interconnect_0:cpu_timer_sw_agent_byteenable -> cpu:timer_sw_agent_byteenable
	wire         mm_interconnect_0_cpu_timer_sw_agent_readdatavalid;        // cpu:timer_sw_agent_readdatavalid -> mm_interconnect_0:cpu_timer_sw_agent_readdatavalid
	wire         mm_interconnect_0_cpu_timer_sw_agent_write;                // mm_interconnect_0:cpu_timer_sw_agent_write -> cpu:timer_sw_agent_write
	wire  [31:0] mm_interconnect_0_cpu_timer_sw_agent_writedata;            // mm_interconnect_0:cpu_timer_sw_agent_writedata -> cpu:timer_sw_agent_writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [15:0] cpu_platform_irq_rx_irq;                                   // irq_mapper:sender_irq -> cpu:platform_irq_rx_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [cpu:reset_reset, data_instruction_ram:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, pio_8bit:reset_n, ram_32bit:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [data_instruction_ram:reset_req, ram_32bit:reset_req, rst_translator:reset_req_in]
	wire         reset_in_out_reset_reset;                                  // reset_in:out_reset -> rst_controller:reset_in0

	sys_clock_in clock_in (
		.in_clk  (clk_clk),              //   input,  width = 1,  in_clk.clk
		.out_clk (clock_in_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	cpu cpu (
		.clk                          (clock_in_out_clk_clk),                               //   input,   width = 1,                 clk.clk
		.reset_reset                  (rst_controller_reset_out_reset),                     //   input,   width = 1,               reset.reset
		.platform_irq_rx_irq          (cpu_platform_irq_rx_irq),                            //   input,  width = 16,     platform_irq_rx.irq
		.instruction_manager_awaddr   (cpu_instruction_manager_awaddr),                     //  output,  width = 32, instruction_manager.awaddr
		.instruction_manager_awsize   (cpu_instruction_manager_awsize),                     //  output,   width = 3,                    .awsize
		.instruction_manager_awprot   (cpu_instruction_manager_awprot),                     //  output,   width = 3,                    .awprot
		.instruction_manager_awvalid  (cpu_instruction_manager_awvalid),                    //  output,   width = 1,                    .awvalid
		.instruction_manager_awready  (cpu_instruction_manager_awready),                    //   input,   width = 1,                    .awready
		.instruction_manager_wdata    (cpu_instruction_manager_wdata),                      //  output,  width = 32,                    .wdata
		.instruction_manager_wstrb    (cpu_instruction_manager_wstrb),                      //  output,   width = 4,                    .wstrb
		.instruction_manager_wlast    (cpu_instruction_manager_wlast),                      //  output,   width = 1,                    .wlast
		.instruction_manager_wvalid   (cpu_instruction_manager_wvalid),                     //  output,   width = 1,                    .wvalid
		.instruction_manager_wready   (cpu_instruction_manager_wready),                     //   input,   width = 1,                    .wready
		.instruction_manager_bresp    (cpu_instruction_manager_bresp),                      //   input,   width = 2,                    .bresp
		.instruction_manager_bvalid   (cpu_instruction_manager_bvalid),                     //   input,   width = 1,                    .bvalid
		.instruction_manager_bready   (cpu_instruction_manager_bready),                     //  output,   width = 1,                    .bready
		.instruction_manager_araddr   (cpu_instruction_manager_araddr),                     //  output,  width = 32,                    .araddr
		.instruction_manager_arsize   (cpu_instruction_manager_arsize),                     //  output,   width = 3,                    .arsize
		.instruction_manager_arprot   (cpu_instruction_manager_arprot),                     //  output,   width = 3,                    .arprot
		.instruction_manager_arvalid  (cpu_instruction_manager_arvalid),                    //  output,   width = 1,                    .arvalid
		.instruction_manager_arready  (cpu_instruction_manager_arready),                    //   input,   width = 1,                    .arready
		.instruction_manager_rdata    (cpu_instruction_manager_rdata),                      //   input,  width = 32,                    .rdata
		.instruction_manager_rresp    (cpu_instruction_manager_rresp),                      //   input,   width = 2,                    .rresp
		.instruction_manager_rvalid   (cpu_instruction_manager_rvalid),                     //   input,   width = 1,                    .rvalid
		.instruction_manager_rready   (cpu_instruction_manager_rready),                     //  output,   width = 1,                    .rready
		.data_manager_awaddr          (cpu_data_manager_awaddr),                            //  output,  width = 32,        data_manager.awaddr
		.data_manager_awsize          (cpu_data_manager_awsize),                            //  output,   width = 3,                    .awsize
		.data_manager_awprot          (cpu_data_manager_awprot),                            //  output,   width = 3,                    .awprot
		.data_manager_awvalid         (cpu_data_manager_awvalid),                           //  output,   width = 1,                    .awvalid
		.data_manager_awready         (cpu_data_manager_awready),                           //   input,   width = 1,                    .awready
		.data_manager_wdata           (cpu_data_manager_wdata),                             //  output,  width = 32,                    .wdata
		.data_manager_wstrb           (cpu_data_manager_wstrb),                             //  output,   width = 4,                    .wstrb
		.data_manager_wlast           (cpu_data_manager_wlast),                             //  output,   width = 1,                    .wlast
		.data_manager_wvalid          (cpu_data_manager_wvalid),                            //  output,   width = 1,                    .wvalid
		.data_manager_wready          (cpu_data_manager_wready),                            //   input,   width = 1,                    .wready
		.data_manager_bresp           (cpu_data_manager_bresp),                             //   input,   width = 2,                    .bresp
		.data_manager_bvalid          (cpu_data_manager_bvalid),                            //   input,   width = 1,                    .bvalid
		.data_manager_bready          (cpu_data_manager_bready),                            //  output,   width = 1,                    .bready
		.data_manager_araddr          (cpu_data_manager_araddr),                            //  output,  width = 32,                    .araddr
		.data_manager_arsize          (cpu_data_manager_arsize),                            //  output,   width = 3,                    .arsize
		.data_manager_arprot          (cpu_data_manager_arprot),                            //  output,   width = 3,                    .arprot
		.data_manager_arvalid         (cpu_data_manager_arvalid),                           //  output,   width = 1,                    .arvalid
		.data_manager_arready         (cpu_data_manager_arready),                           //   input,   width = 1,                    .arready
		.data_manager_rdata           (cpu_data_manager_rdata),                             //   input,  width = 32,                    .rdata
		.data_manager_rresp           (cpu_data_manager_rresp),                             //   input,   width = 2,                    .rresp
		.data_manager_rvalid          (cpu_data_manager_rvalid),                            //   input,   width = 1,                    .rvalid
		.data_manager_rready          (cpu_data_manager_rready),                            //  output,   width = 1,                    .rready
		.timer_sw_agent_write         (mm_interconnect_0_cpu_timer_sw_agent_write),         //   input,   width = 1,      timer_sw_agent.write
		.timer_sw_agent_writedata     (mm_interconnect_0_cpu_timer_sw_agent_writedata),     //   input,  width = 32,                    .writedata
		.timer_sw_agent_byteenable    (mm_interconnect_0_cpu_timer_sw_agent_byteenable),    //   input,   width = 4,                    .byteenable
		.timer_sw_agent_address       (mm_interconnect_0_cpu_timer_sw_agent_address),       //   input,   width = 6,                    .address
		.timer_sw_agent_read          (mm_interconnect_0_cpu_timer_sw_agent_read),          //   input,   width = 1,                    .read
		.timer_sw_agent_readdata      (mm_interconnect_0_cpu_timer_sw_agent_readdata),      //  output,  width = 32,                    .readdata
		.timer_sw_agent_readdatavalid (mm_interconnect_0_cpu_timer_sw_agent_readdatavalid), //  output,   width = 1,                    .readdatavalid
		.dm_agent_write               (mm_interconnect_0_cpu_dm_agent_write),               //   input,   width = 1,            dm_agent.write
		.dm_agent_writedata           (mm_interconnect_0_cpu_dm_agent_writedata),           //   input,  width = 32,                    .writedata
		.dm_agent_address             (mm_interconnect_0_cpu_dm_agent_address),             //   input,  width = 16,                    .address
		.dm_agent_read                (mm_interconnect_0_cpu_dm_agent_read),                //   input,   width = 1,                    .read
		.dm_agent_readdata            (mm_interconnect_0_cpu_dm_agent_readdata),            //  output,  width = 32,                    .readdata
		.dm_agent_readdatavalid       (mm_interconnect_0_cpu_dm_agent_readdatavalid),       //  output,   width = 1,                    .readdatavalid
		.dm_agent_waitrequest         (mm_interconnect_0_cpu_dm_agent_waitrequest)          //  output,   width = 1,                    .waitrequest
	);

	data_instruction_ram data_instruction_ram (
		.clk        (clock_in_out_clk_clk),                                 //   input,   width = 1,   clk1.clk
		.address    (mm_interconnect_0_data_instruction_ram_s1_address),    //   input,  width = 17,     s1.address
		.clken      (mm_interconnect_0_data_instruction_ram_s1_clken),      //   input,   width = 1,       .clken
		.chipselect (mm_interconnect_0_data_instruction_ram_s1_chipselect), //   input,   width = 1,       .chipselect
		.write      (mm_interconnect_0_data_instruction_ram_s1_write),      //   input,   width = 1,       .write
		.readdata   (mm_interconnect_0_data_instruction_ram_s1_readdata),   //  output,  width = 32,       .readdata
		.writedata  (mm_interconnect_0_data_instruction_ram_s1_writedata),  //   input,  width = 32,       .writedata
		.byteenable (mm_interconnect_0_data_instruction_ram_s1_byteenable), //   input,   width = 4,       .byteenable
		.reset      (rst_controller_reset_out_reset),                       //   input,   width = 1, reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                    //   input,   width = 1,       .reset_req
	);

	jtag_uart jtag_uart (
		.clk            (clock_in_out_clk_clk),                                      //   input,   width = 1,               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //   input,   width = 1,             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //   input,   width = 1, avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //   input,   width = 1,                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //   input,   width = 1,                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //  output,  width = 32,                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //   input,   width = 1,                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //   input,  width = 32,                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //  output,   width = 1,                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //  output,   width = 1,               irq.irq
	);

	pio_8bit pio_8bit (
		.clk        (clock_in_out_clk_clk),                     //   input,   width = 1,                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //   input,   width = 1,               reset.reset_n
		.address    (mm_interconnect_0_pio_8bit_s1_address),    //   input,   width = 2,                  s1.address
		.write_n    (~mm_interconnect_0_pio_8bit_s1_write),     //   input,   width = 1,                    .write_n
		.writedata  (mm_interconnect_0_pio_8bit_s1_writedata),  //   input,  width = 32,                    .writedata
		.chipselect (mm_interconnect_0_pio_8bit_s1_chipselect), //   input,   width = 1,                    .chipselect
		.readdata   (mm_interconnect_0_pio_8bit_s1_readdata),   //  output,  width = 32,                    .readdata
		.out_port   (pio_8bit_export)                           //  output,   width = 8, external_connection.export
	);

	ram_32bit ram_32bit (
		.clk        (clock_in_out_clk_clk),                      //   input,   width = 1,   clk1.clk
		.address    (mm_interconnect_0_ram_32bit_s1_address),    //   input,   width = 6,     s1.address
		.clken      (mm_interconnect_0_ram_32bit_s1_clken),      //   input,   width = 1,       .clken
		.chipselect (mm_interconnect_0_ram_32bit_s1_chipselect), //   input,   width = 1,       .chipselect
		.write      (mm_interconnect_0_ram_32bit_s1_write),      //   input,   width = 1,       .write
		.readdata   (mm_interconnect_0_ram_32bit_s1_readdata),   //  output,  width = 32,       .readdata
		.writedata  (mm_interconnect_0_ram_32bit_s1_writedata),  //   input,  width = 32,       .writedata
		.byteenable (mm_interconnect_0_ram_32bit_s1_byteenable), //   input,   width = 4,       .byteenable
		.reset      (rst_controller_reset_out_reset),            //   input,   width = 1, reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)         //   input,   width = 1,       .reset_req
	);

	sys_reset_in reset_in (
		.clk       (clock_in_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset  (reset_reset),              //   input,  width = 1,  in_reset.reset
		.out_reset (reset_in_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	sys_altera_mm_interconnect_1920_5k4ctly mm_interconnect_0 (
		.cpu_data_manager_awaddr                 (cpu_data_manager_awaddr),                                   //   input,  width = 32,                cpu_data_manager.awaddr
		.cpu_data_manager_awsize                 (cpu_data_manager_awsize),                                   //   input,   width = 3,                                .awsize
		.cpu_data_manager_awprot                 (cpu_data_manager_awprot),                                   //   input,   width = 3,                                .awprot
		.cpu_data_manager_awvalid                (cpu_data_manager_awvalid),                                  //   input,   width = 1,                                .awvalid
		.cpu_data_manager_awready                (cpu_data_manager_awready),                                  //  output,   width = 1,                                .awready
		.cpu_data_manager_wdata                  (cpu_data_manager_wdata),                                    //   input,  width = 32,                                .wdata
		.cpu_data_manager_wstrb                  (cpu_data_manager_wstrb),                                    //   input,   width = 4,                                .wstrb
		.cpu_data_manager_wlast                  (cpu_data_manager_wlast),                                    //   input,   width = 1,                                .wlast
		.cpu_data_manager_wvalid                 (cpu_data_manager_wvalid),                                   //   input,   width = 1,                                .wvalid
		.cpu_data_manager_wready                 (cpu_data_manager_wready),                                   //  output,   width = 1,                                .wready
		.cpu_data_manager_bresp                  (cpu_data_manager_bresp),                                    //  output,   width = 2,                                .bresp
		.cpu_data_manager_bvalid                 (cpu_data_manager_bvalid),                                   //  output,   width = 1,                                .bvalid
		.cpu_data_manager_bready                 (cpu_data_manager_bready),                                   //   input,   width = 1,                                .bready
		.cpu_data_manager_araddr                 (cpu_data_manager_araddr),                                   //   input,  width = 32,                                .araddr
		.cpu_data_manager_arsize                 (cpu_data_manager_arsize),                                   //   input,   width = 3,                                .arsize
		.cpu_data_manager_arprot                 (cpu_data_manager_arprot),                                   //   input,   width = 3,                                .arprot
		.cpu_data_manager_arvalid                (cpu_data_manager_arvalid),                                  //   input,   width = 1,                                .arvalid
		.cpu_data_manager_arready                (cpu_data_manager_arready),                                  //  output,   width = 1,                                .arready
		.cpu_data_manager_rdata                  (cpu_data_manager_rdata),                                    //  output,  width = 32,                                .rdata
		.cpu_data_manager_rresp                  (cpu_data_manager_rresp),                                    //  output,   width = 2,                                .rresp
		.cpu_data_manager_rvalid                 (cpu_data_manager_rvalid),                                   //  output,   width = 1,                                .rvalid
		.cpu_data_manager_rready                 (cpu_data_manager_rready),                                   //   input,   width = 1,                                .rready
		.cpu_instruction_manager_awaddr          (cpu_instruction_manager_awaddr),                            //   input,  width = 32,         cpu_instruction_manager.awaddr
		.cpu_instruction_manager_awsize          (cpu_instruction_manager_awsize),                            //   input,   width = 3,                                .awsize
		.cpu_instruction_manager_awprot          (cpu_instruction_manager_awprot),                            //   input,   width = 3,                                .awprot
		.cpu_instruction_manager_awvalid         (cpu_instruction_manager_awvalid),                           //   input,   width = 1,                                .awvalid
		.cpu_instruction_manager_awready         (cpu_instruction_manager_awready),                           //  output,   width = 1,                                .awready
		.cpu_instruction_manager_wdata           (cpu_instruction_manager_wdata),                             //   input,  width = 32,                                .wdata
		.cpu_instruction_manager_wstrb           (cpu_instruction_manager_wstrb),                             //   input,   width = 4,                                .wstrb
		.cpu_instruction_manager_wlast           (cpu_instruction_manager_wlast),                             //   input,   width = 1,                                .wlast
		.cpu_instruction_manager_wvalid          (cpu_instruction_manager_wvalid),                            //   input,   width = 1,                                .wvalid
		.cpu_instruction_manager_wready          (cpu_instruction_manager_wready),                            //  output,   width = 1,                                .wready
		.cpu_instruction_manager_bresp           (cpu_instruction_manager_bresp),                             //  output,   width = 2,                                .bresp
		.cpu_instruction_manager_bvalid          (cpu_instruction_manager_bvalid),                            //  output,   width = 1,                                .bvalid
		.cpu_instruction_manager_bready          (cpu_instruction_manager_bready),                            //   input,   width = 1,                                .bready
		.cpu_instruction_manager_araddr          (cpu_instruction_manager_araddr),                            //   input,  width = 32,                                .araddr
		.cpu_instruction_manager_arsize          (cpu_instruction_manager_arsize),                            //   input,   width = 3,                                .arsize
		.cpu_instruction_manager_arprot          (cpu_instruction_manager_arprot),                            //   input,   width = 3,                                .arprot
		.cpu_instruction_manager_arvalid         (cpu_instruction_manager_arvalid),                           //   input,   width = 1,                                .arvalid
		.cpu_instruction_manager_arready         (cpu_instruction_manager_arready),                           //  output,   width = 1,                                .arready
		.cpu_instruction_manager_rdata           (cpu_instruction_manager_rdata),                             //  output,  width = 32,                                .rdata
		.cpu_instruction_manager_rresp           (cpu_instruction_manager_rresp),                             //  output,   width = 2,                                .rresp
		.cpu_instruction_manager_rvalid          (cpu_instruction_manager_rvalid),                            //  output,   width = 1,                                .rvalid
		.cpu_instruction_manager_rready          (cpu_instruction_manager_rready),                            //   input,   width = 1,                                .rready
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //  output,   width = 1,     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //  output,   width = 1,                                .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //  output,   width = 1,                                .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //   input,  width = 32,                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //  output,  width = 32,                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //   input,   width = 1,                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //  output,   width = 1,                                .chipselect
		.cpu_dm_agent_address                    (mm_interconnect_0_cpu_dm_agent_address),                    //  output,  width = 16,                    cpu_dm_agent.address
		.cpu_dm_agent_write                      (mm_interconnect_0_cpu_dm_agent_write),                      //  output,   width = 1,                                .write
		.cpu_dm_agent_read                       (mm_interconnect_0_cpu_dm_agent_read),                       //  output,   width = 1,                                .read
		.cpu_dm_agent_readdata                   (mm_interconnect_0_cpu_dm_agent_readdata),                   //   input,  width = 32,                                .readdata
		.cpu_dm_agent_writedata                  (mm_interconnect_0_cpu_dm_agent_writedata),                  //  output,  width = 32,                                .writedata
		.cpu_dm_agent_readdatavalid              (mm_interconnect_0_cpu_dm_agent_readdatavalid),              //   input,   width = 1,                                .readdatavalid
		.cpu_dm_agent_waitrequest                (mm_interconnect_0_cpu_dm_agent_waitrequest),                //   input,   width = 1,                                .waitrequest
		.data_instruction_ram_s1_address         (mm_interconnect_0_data_instruction_ram_s1_address),         //  output,  width = 17,         data_instruction_ram_s1.address
		.data_instruction_ram_s1_write           (mm_interconnect_0_data_instruction_ram_s1_write),           //  output,   width = 1,                                .write
		.data_instruction_ram_s1_readdata        (mm_interconnect_0_data_instruction_ram_s1_readdata),        //   input,  width = 32,                                .readdata
		.data_instruction_ram_s1_writedata       (mm_interconnect_0_data_instruction_ram_s1_writedata),       //  output,  width = 32,                                .writedata
		.data_instruction_ram_s1_byteenable      (mm_interconnect_0_data_instruction_ram_s1_byteenable),      //  output,   width = 4,                                .byteenable
		.data_instruction_ram_s1_chipselect      (mm_interconnect_0_data_instruction_ram_s1_chipselect),      //  output,   width = 1,                                .chipselect
		.data_instruction_ram_s1_clken           (mm_interconnect_0_data_instruction_ram_s1_clken),           //  output,   width = 1,                                .clken
		.ram_32bit_s1_address                    (mm_interconnect_0_ram_32bit_s1_address),                    //  output,   width = 6,                    ram_32bit_s1.address
		.ram_32bit_s1_write                      (mm_interconnect_0_ram_32bit_s1_write),                      //  output,   width = 1,                                .write
		.ram_32bit_s1_readdata                   (mm_interconnect_0_ram_32bit_s1_readdata),                   //   input,  width = 32,                                .readdata
		.ram_32bit_s1_writedata                  (mm_interconnect_0_ram_32bit_s1_writedata),                  //  output,  width = 32,                                .writedata
		.ram_32bit_s1_byteenable                 (mm_interconnect_0_ram_32bit_s1_byteenable),                 //  output,   width = 4,                                .byteenable
		.ram_32bit_s1_chipselect                 (mm_interconnect_0_ram_32bit_s1_chipselect),                 //  output,   width = 1,                                .chipselect
		.ram_32bit_s1_clken                      (mm_interconnect_0_ram_32bit_s1_clken),                      //  output,   width = 1,                                .clken
		.pio_8bit_s1_address                     (mm_interconnect_0_pio_8bit_s1_address),                     //  output,   width = 2,                     pio_8bit_s1.address
		.pio_8bit_s1_write                       (mm_interconnect_0_pio_8bit_s1_write),                       //  output,   width = 1,                                .write
		.pio_8bit_s1_readdata                    (mm_interconnect_0_pio_8bit_s1_readdata),                    //   input,  width = 32,                                .readdata
		.pio_8bit_s1_writedata                   (mm_interconnect_0_pio_8bit_s1_writedata),                   //  output,  width = 32,                                .writedata
		.pio_8bit_s1_chipselect                  (mm_interconnect_0_pio_8bit_s1_chipselect),                  //  output,   width = 1,                                .chipselect
		.cpu_timer_sw_agent_address              (mm_interconnect_0_cpu_timer_sw_agent_address),              //  output,   width = 6,              cpu_timer_sw_agent.address
		.cpu_timer_sw_agent_write                (mm_interconnect_0_cpu_timer_sw_agent_write),                //  output,   width = 1,                                .write
		.cpu_timer_sw_agent_read                 (mm_interconnect_0_cpu_timer_sw_agent_read),                 //  output,   width = 1,                                .read
		.cpu_timer_sw_agent_readdata             (mm_interconnect_0_cpu_timer_sw_agent_readdata),             //   input,  width = 32,                                .readdata
		.cpu_timer_sw_agent_writedata            (mm_interconnect_0_cpu_timer_sw_agent_writedata),            //  output,  width = 32,                                .writedata
		.cpu_timer_sw_agent_byteenable           (mm_interconnect_0_cpu_timer_sw_agent_byteenable),           //  output,   width = 4,                                .byteenable
		.cpu_timer_sw_agent_readdatavalid        (mm_interconnect_0_cpu_timer_sw_agent_readdatavalid),        //   input,   width = 1,                                .readdatavalid
		.cpu_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            //   input,   width = 1, cpu_reset_reset_bridge_in_reset.reset
		.clock_in_out_clk_clk                    (clock_in_out_clk_clk)                                       //   input,   width = 1,                clock_in_out_clk.clk
	);

	sys_altera_irq_mapper_1920_jj7diii irq_mapper (
		.clk           (clock_in_out_clk_clk),           //   input,   width = 1,       clk.clk
		.reset         (rst_controller_reset_out_reset), //   input,   width = 1, clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       //   input,   width = 1, receiver0.irq
		.sender_irq    (cpu_platform_irq_rx_irq)         //  output,  width = 16,    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_in_out_reset_reset),           //   input,  width = 1, reset_in0.reset
		.clk            (clock_in_out_clk_clk),               //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
